//	setup file time 2018/2/6
//	author <ross1206vii@gmail.com>



module select_16
(
	in,
	sel,
	out
);


input[15:0] in;
input[3:0] sel;
output out;



always @(*)
begin
//	case(sel)
//		4'b0000:
//			out = in[0];
	
	
//	endcase
end



endmodule

